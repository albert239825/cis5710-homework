/* INSERT NAME AND PENNKEY HERE */

`timescale 1ns / 1ns

// quotient = dividend / divisor

module DividerUnsigned (
    input  wire [31:0] i_dividend,
    input  wire [31:0] i_divisor,
    output wire [31:0] o_remainder,
    output wire [31:0] o_quotient
);

    // TODO: your code here

endmodule


module DividerOneIter (
    input  wire [31:0] i_dividend,
    input  wire [31:0] i_divisor,
    input  wire [31:0] i_remainder,
    input  wire [31:0] i_quotient,
    output logic [31:0] o_dividend,
    output logic [31:0] o_remainder,
    output logic [31:0] o_quotient
);
  /*
    for (int i = 0; i < 32; i++) {
        remainder = (remainder << 1) | ((dividend >> 31) & 0x1);
        if (remainder < divisor) {
            quotient = (quotient << 1);
        } else {
            quotient = (quotient << 1) | 0x1;
            remainder = remainder - divisor;
        }
        dividend = dividend << 1;
    }
    */

    // TODO: your code here

    logic [31:0] rem_shift;

    always_comb begin
        rem_shift = i_remainder << 1 | {31'b0, i_dividend[31]};
        if (rem_shift < i_divisor) begin
            o_quotient = i_quotient << 1;
            o_remainder = rem_shift;
        end else begin
            o_quotient = {i_quotient[31:1], 1'b1};
            o_remainder = rem_shift - i_divisor;
        end
        o_dividend = {i_dividend[31:1], 1'b0};
    end

endmodule
